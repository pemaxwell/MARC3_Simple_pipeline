reset_vector_inst : reset_vector PORT MAP (
		result	 => result_sig
	);
