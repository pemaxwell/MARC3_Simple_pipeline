--------------------------------------------------------------------------------------		
--		File:  CPU_chip.vhd
--
--		Created by: MAJ Paul Maxwell
--
--		Date Created:  4 Sep 03
--
--		Modified by:  LTC Paul Maxwell
--
--		Date Last Modified:  5 Jun 2012
--
--		Version:  2.0
--
-- 	Description:  This file provides the top-level design for the EE375 MARC2 
--			processor.  Using the constraints file provided and this code, the user can
--			insert a cadet's MARC2 source code into this project (replacing my cpu_marc1
--			and its dependent files) and implement this processor in hardware.  This 
--			solution is designed for an Altera Cyclone IVE chip on an 
--			Terasic DE2-115 Education and Development Board.  
--
-------------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity CPU_chip is
    Port ( 	clk : in std_logic;   										-- CPU clock
				reset : in std_logic;			 							-- Key0
				run : in std_logic;			 								-- SW17 
				reg_select : in std_LOGIC_VECTOR(2 downto 0);		-- SW2-SW0 (LSb), select lines for register output
				LCD_RS, LCD_E, LCD_ON, LCD_RW, RESET_LED, SEC_LED : out std_LOGIC; --lcd control signals
				lcd_data : INOUT	STD_LOGIC_VECTOR(7 DOWNTO 0)  	-- data lines to lcd displayReg
			);
end CPU_chip;

architecture Behavioral of CPU_chip is

component CPU_MARC1 is
    port (
		clk: IN std_logic;					-- system clock
		mem_rd : OUT std_logic;				-- memory read control
		mem_wr : OUT std_logic;				-- memory write control  
		mem_cs : OUT std_logic;				-- memory chip select
		address: INOUT std_logic_vector(15 downto 0); -- system addr bus
		data: INOUT std_logic_vector(15 downto 0);  -- system data bus
		R1out,R2out,R3out,R4out,R5out,R6out,R7out : out std_logic_vector(15 downto 0);
		run : IN std_logic;   				-- external run signal
		rst: IN  std_logic	  				-- external reset signal
     ); 
end component;

--  The following RAM and ROM are generated by the Coregen tool.  They are created as
--	 single port block memory units which are clocked on the falling edge in order to 
--	 remove some timing conflicts.

component systemram 
	PORT
	(
		address	: IN STD_LOGIC_VECTOR (10 DOWNTO 0);
		clock		: IN STD_LOGIC  := '1';
		data		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		wren		: IN STD_LOGIC ;
		q			: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
END component;


component systemrom 
	PORT
	(
		address	: IN STD_LOGIC_VECTOR (9 DOWNTO 0);
		clock		: IN STD_LOGIC  := '1';
		q			: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
END component;

component DE2_CLOCK 
	PORT(
			reset, clk_50Mhz	: IN	STD_LOGIC;
			LCD_RS, LCD_E, LCD_ON, RESET_LED	: OUT	STD_LOGIC;
			LCD_RW				: BUFFER STD_LOGIC;
			display_data		: IN std_LOGIC_VECTOR(15 downto 0);
			DATA_BUS				: INOUT	STD_LOGIC_VECTOR(7 DOWNTO 0)
		  );
END component;

signal Addr_bus, Data_bus, data_bus_temp, data_out1,data_out2, dummy : std_logic_vector(15 downto 0);  --TEST_IT, B_bus, PC,
signal mem_rd, mem_wr, mem_cs, mem_cs_ram, mem_cs_rom, divclkout, runSp, rstSP : std_logic;
signal R1out,R2out,R3out,R4out,R5out,R6out,R7out,DisplayReg : std_logic_vector(15 downto 0);
signal AddrOut, DataOut, RegOut, InfoOut : std_logic_vector(6 downto 0);
signal AddrHex, DataHex, RegHex, RegSel : std_logic_vector(3 downto 0);
signal display_buf : std_logic_vector(15 downto 0);
signal system_clock, memory_clk : std_LOGIC;			--added 21 Nov 12 to deal with double registered memory


begin

runSP <= run;						--switch set to exterior of board = off (don't run); 
rstSP <= reset;					--changed to reflect that pushbutton outputs '1' when button isn't pushed 13 Nov 12
SEC_LED <= '1';
memory_clk <= clk;

sys_clk_divider: process (clk, reset)
begin
	if (reset = '0') then system_clock <= '1'; 
	elsif (rising_edge(clk) and clk = '1')then
		system_clock <= not system_clock;
	end if;
end process;


mem_cs_rom <= '1' when ((mem_cs='0')and(mem_rd='0')and(addr_bus(12 downto 10)="000")) else
				  '0';

mem_cs_ram <= '1' when ((mem_cs='0')and(mem_rd='0')and((addr_bus(12 downto 10)="001")or
					(addr_bus(12 downto 10)="100")or(addr_bus(12 downto 10)="010")or
					(addr_bus(12 downto 10)="011"))) else
				  '0';

data_bus_temp <= data_out1 when mem_cs_ram = '1' else
				     data_out2 when mem_cs_rom = '1' else
					  "ZZZZZZZZZZZZZZZZ";
					  
displayReg <= R1out when reg_select = "001" else
					R2out when reg_select = "010" else
					R3out when reg_select = "011" else
					R4out when reg_select = "100" else
					R5out when reg_select = "101" else	
					R6out when reg_select = "110" else
					R7out when reg_select = "111" else
					display_buf;

Ram1 : systemram
		port map (address => addr_bus(10 downto 0), clock => memory_clk, data => data_bus_temp,
			q => data_out1, wren => mem_wr);

ProgMem : systemrom
		port map (address => addr_bus(9 downto 0), clock => memory_clk, q => data_out2);

CPU: CPU_MARC1 port map(system_clock, mem_rd, mem_wr,mem_cs, addr_bus,	data_bus_temp,R1out,R2out,
			R3out,R4out,R5out,R6out,R7out,runSP,rstSP); 	
			
lcd_out:  DE2_CLOCK port map( reset, clk, LCD_RS, LCD_E, LCD_ON, RESET_LED, lcd_rw, displayReg, lcd_data);
		  
process (clk, addr_bus)
begin
	if (rising_edge(clk) and addr_bus = X"0800")then
		display_buf <= data_bus_temp;
	end if;
end process;

end Behavioral;
