bit16_2_to_1_mux_inst : bit16_2_to_1_mux PORT MAP (
		data0x	 => data0x_sig,
		data1x	 => data1x_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
