PC_displ_adder_inst : PC_displ_adder PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);
