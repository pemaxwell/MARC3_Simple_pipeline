constant0_inst : constant0 PORT MAP (
		result	 => result_sig
	);
