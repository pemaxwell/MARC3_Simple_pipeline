PC_adder_inst : PC_adder PORT MAP (
		dataa	 => dataa_sig,
		result	 => result_sig
	);
