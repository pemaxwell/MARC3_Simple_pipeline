bit_1_inst : bit_1 PORT MAP (
		result	 => result_sig
	);
