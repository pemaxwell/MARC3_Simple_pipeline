constant1_inst : constant1 PORT MAP (
		result	 => result_sig
	);
