sp_sub_inst : sp_sub PORT MAP (
		dataa	 => dataa_sig,
		result	 => result_sig
	);
